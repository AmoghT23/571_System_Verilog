module testDays();
  reg [4:0]m;
  reg LY;
  wire d27, d28;
  
  DaysDetector d(m, LY, d27, d28);
  
  initial 
    begin
      
      $dumpfile("dump.vcd");
      $dumpvars(1);
      
      #10 LY = 1'bx;
      #10 m=5'b00000;
      #10 m=5'b00001;
      #10 m=5'b00010;
      #10 m=5'b00011;
      #10 m=5'b00100;
      #10 m=5'b00101;
      #10 m=5'b00110;
      #10 m=5'b00111;
      #10 m=5'b01000;
      #10 m=5'b01001;
      #10 m=5'b01010;
      #10 m=5'b01011;
      #10 m=5'b01100;
      #10 m=5'b01101;
      #10 m=5'b01110;
      #10 m=5'b01111;
      #10 m=5'b10000;
      #10 m=5'b10001;
      #10 m=5'b10010;
      #10 m=5'b10011;
      #10 m=5'b10100;
      #10 m=5'b10101;
      #10 m=5'b10110;
      #10 m=5'b10111;
     	#10 LY = 1'b0;
      	#10 LY = 1'b1;
      	#10 LY = 1'bx;
      #10 m=5'b11000;
      #10 m=5'b11001;
      #10 m=5'b11010;
      #10 m=5'b11011;
      #10 m=5'b11100;
      #10 m=5'b11101;
      #10 m=5'b11110;
      #10 m=5'b11111;
      
      $monitor("The binary Value is= %b, d27 = %b",LY,d27);
    end
endmodule
